* C:\Users\mamat\OneDrive\Documents\Final_project_files\Device_Modelling\2N5401\BJT_CB_config_input_char_2N5401\BJT_CB_config_input_char_2N5401.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/17/25 11:15:48

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v1  GND vcb DC		
R1  vcb Net-_Q1-Pad1_ 1k		
R2  Net-_Q1-Pad3_ Net-_R2-Pad2_ 1k		
U_ic1  ie Net-_R2-Pad2_ plot_i2		
v2  ie GND DC		
Q1  Net-_Q1-Pad1_ GND Net-_Q1-Pad3_ eSim_PNP		

.end
