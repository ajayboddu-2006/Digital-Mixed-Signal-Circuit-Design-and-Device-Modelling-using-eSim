* C:\Users\mamat\eSim-Workspace\SN74100_Bistable_Latch\SN74100_Bistable_Latch.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/02/25 12:09:26

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U4  Net-_U4-Pad1_ OUT dac_bridge_1		
U3  D EN Net-_U3-Pad3_ Net-_U3-Pad4_ adc_bridge_2		
v1  D GND pulse		
v2  EN GND pulse		
U1  D plot_v1		
U2  EN plot_v1		
U5  OUT plot_v1		
X1  ? ? ? ? ? ? GND ? ? ? ? ? ? ? ? ? ? ? ? Net-_U4-Pad1_ Net-_U3-Pad3_ ? Net-_U3-Pad4_ Net-_X1-Pad24_ SN74100		
v3  Net-_X1-Pad24_ GND 5		

.end
