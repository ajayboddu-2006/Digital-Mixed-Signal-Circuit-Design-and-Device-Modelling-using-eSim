* C:\Users\mamat\eSim-Workspace\BJT_CE_config_input_char_ZTX1048A\BJT_CE_config_input_char_ZTX1048A.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/13/25 15:27:49

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U_ic1  ib Net-_R1-Pad1_ plot_i2		
Q1  Net-_Q1-Pad1_ Net-_Q1-Pad2_ GND eSim_NPN		
v2  ib GND DC		
R2  vce Net-_Q1-Pad1_ 1k		
R1  Net-_R1-Pad1_ Net-_Q1-Pad2_ 1k		
v1  vce GND DC		

.end
