* C:\Users\mamat\OneDrive\Desktop\Ajay_eSim\Final_project_files\Device_Modelling\2N5401\BJT_CE_config\BJT_CE_config.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/13/25 19:14:27

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v1  GND vce DC		
R1  vce Net-_Q1-Pad1_ 1k		
R2  Net-_Q1-Pad2_ Net-_R2-Pad2_ 1k		
U_ic1  Net-_R2-Pad2_ ib plot_i2		
Q1  Net-_Q1-Pad1_ Net-_Q1-Pad2_ GND eSim_PNP		
v2  GND ib DC		

.end
