* C:\Users\mamat\OneDrive\Documents\Final_project_files\Device_Modelling\2N5401\BJT_CB_config_output_cha_2N5401\BJT_CB_config_output_cha_2N5401.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/17/25 11:20:21

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v1  GND vcb DC		
R1  Net-_R1-Pad1_ Net-_Q1-Pad1_ 1k		
R2  Net-_Q1-Pad3_ ie 1k		
U_ic1  Net-_R1-Pad1_ vcb plot_i2		
I1  ie GND dc		
Q1  Net-_Q1-Pad1_ GND Net-_Q1-Pad3_ eSim_PNP		

.end
