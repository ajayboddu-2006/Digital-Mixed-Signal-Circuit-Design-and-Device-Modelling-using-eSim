* C:\Users\mamat\OneDrive\Documents\Final_project_files\Device_Modelling\PMEG2005EB\Diode_char_PMEG2005EB\Diode_char_PMEG2005EB.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/24/25 15:33:34

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  out Net-_R1-Pad1_ plot_i2		
D1  out in eSim_Diode		
v1  in GND DC		
R1  Net-_R1-Pad1_ GND 1k		

.end
