* C:\Users\Chaithu\FOSSEE\eSim\library\SubcircuitLibrary\ajay\ajay.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 6/1/2025 10:40:05 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U5  Net-_U1-Pad3_ Net-_U3-Pad2_ d_inverter		
U7  Net-_U1-Pad3_ Net-_U1-Pad2_ Net-_U7-Pad3_ d_and		
U3  Net-_U1-Pad2_ Net-_U3-Pad2_ Net-_U2-Pad2_ d_and		
U2  Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U1-Pad1_ d_nor		
U4  Net-_U4-Pad1_ Net-_U2-Pad1_ d_buffer		
U6  Net-_U1-Pad1_ Net-_U6-Pad2_ d_buffer		
U8  Net-_U7-Pad3_ Net-_U6-Pad2_ Net-_U4-Pad1_ d_nor		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ PORT		

.end
